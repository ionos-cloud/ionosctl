module github.com/ionos-cloud/ionosctl

go 1.18

require (
	github.com/cheggaaa/pb/v3 v3.1.0
	github.com/fatih/color v1.13.0
	github.com/fatih/structs v1.1.0
	github.com/golang/mock v1.6.0
	github.com/google/uuid v1.3.0
	github.com/ionos-cloud/sdk-go-auth v1.0.5
	github.com/ionos-cloud/sdk-go-dbaas-postgres v1.0.4
	github.com/ionos-cloud/sdk-go/v6 v6.1.3
	github.com/mitchellh/go-homedir v1.1.0
	github.com/spf13/cobra v1.5.0
	github.com/spf13/pflag v1.0.5
	github.com/spf13/viper v1.13.0
	github.com/stretchr/testify v1.8.0
	github.com/webguerilla/ftps v0.0.0-20180713194618-60e520f5feed
	go.uber.org/multierr v1.8.0
	golang.org/x/crypto v0.0.0-20220919173607-35f4265a4bc0
	golang.org/x/exp v0.0.0-20220921164117-439092de6870
	golang.org/x/term v0.0.0-20220919170432-7a66f970e087
)

require (
	github.com/VividCortex/ewma v1.2.0 // indirect
	github.com/davecgh/go-spew v1.1.1 // indirect
	github.com/fsnotify/fsnotify v1.5.4 // indirect
	github.com/golang/protobuf v1.5.2 // indirect
	github.com/hashicorp/hcl v1.0.0 // indirect
	github.com/inconshreveable/mousetrap v1.0.1 // indirect
	github.com/magiconair/properties v1.8.6 // indirect
	github.com/mattn/go-colorable v0.1.13 // indirect
	github.com/mattn/go-isatty v0.0.16 // indirect
	github.com/mattn/go-runewidth v0.0.14 // indirect
	github.com/mitchellh/mapstructure v1.5.0 // indirect
	github.com/pelletier/go-toml v1.9.5 // indirect
	github.com/pelletier/go-toml/v2 v2.0.5 // indirect
	github.com/pmezard/go-difflib v1.0.0 // indirect
	github.com/rivo/uniseg v0.4.2 // indirect
	github.com/spf13/afero v1.9.2 // indirect
	github.com/spf13/cast v1.5.0 // indirect
	github.com/spf13/jwalterweatherman v1.1.0 // indirect
	github.com/subosito/gotenv v1.4.1 // indirect
	go.uber.org/atomic v1.10.0 // indirect
	golang.org/x/net v0.0.0-20220921203646-d300de134e69 // indirect
	golang.org/x/oauth2 v0.0.0-20220909003341-f21342109be1 // indirect
	golang.org/x/sys v0.0.0-20220919091848-fb04ddd9f9c8 // indirect
	golang.org/x/text v0.3.7 // indirect
	google.golang.org/appengine v1.6.7 // indirect
	google.golang.org/protobuf v1.28.1 // indirect
	gopkg.in/ini.v1 v1.67.0 // indirect
	gopkg.in/yaml.v2 v2.4.0 // indirect
	gopkg.in/yaml.v3 v3.0.1 // indirect
)
